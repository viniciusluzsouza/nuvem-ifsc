library ieee;
use ieee.std_logic_1164.all;
entity shift3mode is
   port(
      a: in std_logic_vector(63 downto 0);
      lar: in std_logic_vector(1 downto 0);
      amt: in std_logic_vector(5 downto 0);
      y: out std_logic_vector(63 downto 0)
   );
end shift3mode ;

--=============================
-- Listing 7.13 barrel shifter
--=============================
architecture direct_arch of shift3mode is
   signal logic_result, arith_result, rot_result:
      std_logic_vector(63 downto 0);
begin
   with amt select
       rot_result<=
          a                                when "000000",
          a(0) & a(63 downto 1)            when "000001",
          a(1 downto 0) & a(63 downto 2)   when "000010",
          a(2 downto 0) & a(63 downto 3)   when "000011",
          a(3 downto 0) & a(63 downto 4)   when "000100",
          a(4 downto 0) & a(63 downto 5)   when "000101",
          a(5 downto 0) & a(63 downto 6)   when "000110",
          a(6 downto 0) & a(63 downto 7)   when "000111",
			 a(7 downto 0) & a(63 downto 8)   when "001000",
          a(8 downto 0) & a(63 downto 9)   when "001001",
          a(9 downto 0) & a(63 downto 10)  when "001010",
          a(10 downto 0) & a(63 downto 11) when "001011",
          a(11 downto 0) & a(63 downto 12) when "001100",
          a(12 downto 0) & a(63 downto 13) when "001101",
          a(13 downto 0) & a(63 downto 14) when "001110",
          a(14 downto 0) & a(63 downto 15) when "001111",
          a(15 downto 0) & a(63 downto 16) when "010000",
          a(16 downto 0) & a(63 downto 17) when "010001",
          a(17 downto 0) & a(63 downto 18) when "010010",
          a(18 downto 0) & a(63 downto 19) when "010011",
          a(19 downto 0) & a(63 downto 20) when "010100",
          a(20 downto 0) & a(63 downto 21) when "010101",
          a(21 downto 0) & a(63 downto 22) when "010110",
          a(22 downto 0) & a(63 downto 23) when "010111",
			 a(23 downto 0) & a(63 downto 24) when "011000",
          a(24 downto 0) & a(63 downto 25) when "011001",
          a(25 downto 0) & a(63 downto 26) when "011010",
          a(26 downto 0) & a(63 downto 27) when "011011",
          a(27 downto 0) & a(63 downto 28) when "011100",
          a(28 downto 0) & a(63 downto 29) when "011101",
          a(29 downto 0) & a(63 downto 30) when "011110",
          a(30 downto 0) & a(63 downto 31) when "011111",
          a(31 downto 0) & a(63 downto 32) when "100000",
          a(32 downto 0) & a(63 downto 33) when "100001",
          a(33 downto 0) & a(63 downto 34) when "100010",
          a(34 downto 0) & a(63 downto 35) when "100011",
          a(35 downto 0) & a(63 downto 36) when "100100",
          a(36 downto 0) & a(63 downto 37) when "100101",
          a(37 downto 0) & a(63 downto 38) when "100110",
          a(38 downto 0) & a(63 downto 39) when "100111",
			 a(39 downto 0) & a(63 downto 40) when "101000",
          a(40 downto 0) & a(63 downto 41) when "101001",
          a(41 downto 0) & a(63 downto 42) when "101010",
          a(42 downto 0) & a(63 downto 43) when "101011",
          a(43 downto 0) & a(63 downto 44) when "101100",
          a(44 downto 0) & a(63 downto 45) when "101101",
          a(45 downto 0) & a(63 downto 46) when "101110",
          a(46 downto 0) & a(63 downto 47) when "101111",
          a(47 downto 0) & a(63 downto 48) when "110000",
          a(48 downto 0) & a(63 downto 49) when "110001",
          a(49 downto 0) & a(63 downto 50) when "110010",
          a(50 downto 0) & a(63 downto 51) when "110011",
          a(51 downto 0) & a(63 downto 52) when "110100",
          a(52 downto 0) & a(63 downto 53) when "110101",
          a(53 downto 0) & a(63 downto 54) when "110110",
          a(54 downto 0) & a(63 downto 55) when "110111",
			 a(55 downto 0) & a(63 downto 56) when "111000",
          a(56 downto 0) & a(63 downto 57) when "111001",
          a(57 downto 0) & a(63 downto 58) when "111010",
          a(58 downto 0) & a(63 downto 59) when "111011",
          a(59 downto 0) & a(63 downto 60) when "111100",
          a(60 downto 0) & a(63 downto 61) when "111101",
          a(61 downto 0) & a(63 downto 62) when "111110",
          a(62 downto 0) & a(63) when others; -- "111111"

   with amt select
      logic_result<=
          a                    when "000000",
          "0" & a(63 downto 1)  when "000001",
          "00" & a(63 downto 2)  when "000010",
          "000" & a(63 downto 3)  when "000011",
          "0000" & a(63 downto 4)  when "000100",
          "00000" & a(63 downto 5)  when "000101",
          "000000" & a(63 downto 6)  when "000110",
          "0000000" & a(63 downto 7)  when "000111",
			 "00000000" & a(63 downto 8)  when "001000",
          "000000000" & a(63 downto 9)  when "001001",
          "0000000000" & a(63 downto 10) when "001010",
          "00000000000" & a(63 downto 11) when "001011",
          "000000000000" & a(63 downto 12) when "001100",
          "0000000000000" & a(63 downto 13) when "001101",
          "00000000000000" & a(63 downto 14) when "001110",
          "000000000000000" & a(63 downto 15) when "001111",
          "0000000000000000" & a(63 downto 16) when "010000",
          "00000000000000000" & a(63 downto 17) when "010001",
          "000000000000000000" & a(63 downto 18) when "010010",
          "0000000000000000000" & a(63 downto 19) when "010011",
          "00000000000000000000" & a(63 downto 20) when "010100",
          "000000000000000000000" & a(63 downto 21) when "010101",
          "0000000000000000000000" & a(63 downto 22) when "010110",
          "00000000000000000000000" & a(63 downto 23) when "010111",
			 "000000000000000000000000" & a(63 downto 24) when "011000",
          "0000000000000000000000000" & a(63 downto 25) when "011001",
          "00000000000000000000000000" & a(63 downto 26) when "011010",
          "000000000000000000000000000" & a(63 downto 27) when "011011",
          "0000000000000000000000000000" & a(63 downto 28) when "011100",
          "00000000000000000000000000000" & a(63 downto 29) when "011101",
          "000000000000000000000000000000" & a(63 downto 30) when "011110",
          "0000000000000000000000000000000" & a(63 downto 31) when "011111",
          "00000000000000000000000000000000" & a(63 downto 32) when "100000",
          "000000000000000000000000000000000" & a(63 downto 33) when "100001",
          "0000000000000000000000000000000000" & a(63 downto 34) when "100010",
          "00000000000000000000000000000000000" & a(63 downto 35) when "100011",
          "000000000000000000000000000000000000" & a(63 downto 36) when "100100",
          "0000000000000000000000000000000000000" & a(63 downto 37) when "100101",
          "00000000000000000000000000000000000000" & a(63 downto 38) when "100110",
          "000000000000000000000000000000000000000" & a(63 downto 39) when "100111",
			 "0000000000000000000000000000000000000000" & a(63 downto 40) when "101000",
          "00000000000000000000000000000000000000000" & a(63 downto 41) when "101001",
          "000000000000000000000000000000000000000000" & a(63 downto 42) when "101010",
          "0000000000000000000000000000000000000000000" & a(63 downto 43) when "101011",
          "00000000000000000000000000000000000000000000" & a(63 downto 44) when "101100",
          "000000000000000000000000000000000000000000000" & a(63 downto 45) when "101101",
          "0000000000000000000000000000000000000000000000" & a(63 downto 46) when "101110",
          "00000000000000000000000000000000000000000000000" & a(63 downto 47) when "101111",
          "000000000000000000000000000000000000000000000000" & a(63 downto 48) when "110000",
          "0000000000000000000000000000000000000000000000000" & a(63 downto 49) when "110001",
          "00000000000000000000000000000000000000000000000000" & a(63 downto 50) when "110010",
          "000000000000000000000000000000000000000000000000000" & a(63 downto 51) when "110011",
          "0000000000000000000000000000000000000000000000000000" & a(63 downto 52) when "110100",
          "00000000000000000000000000000000000000000000000000000" & a(63 downto 53) when "110101",
          "000000000000000000000000000000000000000000000000000000" & a(63 downto 54) when "110110",
          "0000000000000000000000000000000000000000000000000000000" & a(63 downto 55) when "110111",
			 "00000000000000000000000000000000000000000000000000000000" & a(63 downto 56) when "111000",
          "000000000000000000000000000000000000000000000000000000000" & a(63 downto 57) when "111001",
          "0000000000000000000000000000000000000000000000000000000000" & a(63 downto 58) when "111010",
          "00000000000000000000000000000000000000000000000000000000000" & a(63 downto 59) when "111011",
          "000000000000000000000000000000000000000000000000000000000000" & a(63 downto 60) when "111100",
          "0000000000000000000000000000000000000000000000000000000000000" & a(63 downto 61) when "111101",
          "00000000000000000000000000000000000000000000000000000000000000" & a(63 downto 62) when "111110",
          "000000000000000000000000000000000000000000000000000000000000000" & a(63) when others; -- "111111"

   with amt select
      arith_result<=
         a               when "000000",
			a(63)& a(63 downto 1) when "000001",
			a(63)&a(63)& a(63 downto 2) when "000010",
			a(63)&a(63)&a(63)& a(63 downto 3) when "000011",
			a(63)&a(63)&a(63)&a(63)& a(63 downto 4) when "000100",
			a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 5) when "000101",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 6) when "000110",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 7) when "000111",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 8) when "001000",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 9) when "001001",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 10) when "001010",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 11) when "001011",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 12) when "001100",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 13) when "001101",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 14) when "001110",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 15) when "001111",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 16) when "010000",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 17) when "010001",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 18) when "010010",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 19) when "010011",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 20) when "010100",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 21) when "010101",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 22) when "010110",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 23) when "010111",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 24) when "011000",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 25) when "011001",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 26) when "011010",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 27) when "011011",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 28) when "011100",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 29) when "011101",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 30) when "011110",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 31) when "011111",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 32) when "100000",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 33) when "100001",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 34) when "100010",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 35) when "100011",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 36) when "100100",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 37) when "100101",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 38) when "100110",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 39) when "100111",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 40) when "101000",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 41) when "101001",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 42) when "101010",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 43) when "101011",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 44) when "101100",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 45) when "101101",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 46) when "101110",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 47) when "101111",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 48) when "110000",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 49) when "110001",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 50) when "110010",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 51) when "110011",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 52) when "110100",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 53) when "110101",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 54) when "110110",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 55) when "110111",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 56) when "111000",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 57) when "111001",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 58) when "111010",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 59) when "111011",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 60) when "111100",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 61) when "111101",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63 downto 62) when "111110",
			a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)&a(63)& a(63) when others; -- "111111"
   with lar select
      y <= logic_result when "00",
           arith_result when "01",
           rot_result   when others;
end direct_arch;