    Mac OS X            	   2   �                                           ATTR         �                     �     com.apple.lastuseddate#PS           com.macromates.selectionRange           com.macromates.visibleIndex  ���Z    _�    10