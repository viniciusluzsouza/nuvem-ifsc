    Mac OS X            	   2   �                                           ATTR         �                     �     com.apple.lastuseddate#PS           com.macromates.selectionRange      	     com.macromates.visibleIndex  2��Z    C�    17:22712